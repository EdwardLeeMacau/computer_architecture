module ALU_Control
(

);

endmodule
