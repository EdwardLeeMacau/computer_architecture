module Branch_Predictor
(
    output              predict_o
);

assign predict_o = 1'b0;

endmodule