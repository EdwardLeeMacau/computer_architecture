module Control
(

);

endmodule
