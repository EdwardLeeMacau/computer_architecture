module MUX32
(

);

endmodule
