module ALU
(

);

endmodule