module Sign_Extend
(

);

endmodule
