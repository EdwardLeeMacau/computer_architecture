module Adder
(

);

endmodule
